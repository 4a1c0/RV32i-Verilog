@00000000
13 01 01 FE 23 2E 81 00 13 04 01 02 23 26 04 FE 
93 07 40 01 23 24 F4 FE 23 26 04 FE 6F 00 C0 01 
83 27 84 FE 03 27 C4 FE 23 A0 E7 00 83 27 C4 FE 
93 87 17 00 23 26 F4 FE 03 27 C4 FE 93 07 F0 01 
E3 D0 E7 FE 83 27 84 FE 13 07 F0 1F 23 A0 E7 00 
93 07 00 00 13 85 07 00 03 24 C1 01 13 01 01 02 
67 80 00 00 
